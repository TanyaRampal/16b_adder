/home/t3rampal/ECE637/cadence/proj2_1bit_fulladder/lvs/netlist